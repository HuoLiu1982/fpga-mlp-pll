`timescale 1ns/1ps

module dblcordicpll_top (
    // ʱ�Ӻ͸�λ
    input  wire         clk,           // ϵͳʱ��
    input  wire         reset_n,       // �첽��λ���͵�ƽ��Ч
    input  wire         enable_posedge,        // AD����ʱ�ӵ������أ�������Ч�źţ�
    
    // �����ź�
    input  wire signed [15:0] signal_in,  // �����ź�
    input  wire          r_error_jump,        // ���ͻ���־ 
    // ����ź�
    output wire [15:0]  phase_error,   // ��λ���ȶ�ֵ2**15
    output wire [31:0]  output_phase,   // �����λ
    output wire         pll_done
    
);

    // ��������
    parameter IW = 16;      // ����λ��
    parameter PW = 32;      // ��λλ��  
    parameter OW = 16;      // ���λ��
    
    // ����ϵ������ - ��3��14
    localparam GAIN_3  = 5'd3;     // ����3
    localparam GAIN_4  = 5'd4;     // ����4
    localparam GAIN_5  = 5'd5;     // ����5
    localparam GAIN_6  = 5'd6;     // ����6
    localparam GAIN_7  = 5'd7;     // ����7
    localparam GAIN_8  = 5'd8;     // ����8
    localparam GAIN_9  = 5'd9;     // ����9
    localparam GAIN_10 = 5'd10;    // ����10
    localparam GAIN_11 = 5'd11;    // ����11
    localparam GAIN_12 = 5'd12;    // ����12
    localparam GAIN_13 = 5'd13;    // ����13
    localparam GAIN_14 = 5'd14;    // ����14
    
    // ����ʱ�䱶������ - ��������Ҫ�����
    localparam DUL_3_TO_4   = 32'd3;    // 3->4: 1��
    localparam DUL_4_TO_5   = 32'd3;    // 4->5: 1��
    localparam DUL_5_TO_6   = 32'd3;    // 5->6: 1��
    localparam DUL_6_TO_7   = 32'd3;    // 6->7: 3��
    localparam DUL_7_TO_8   = 32'd3;    // 7->8: 3��
    localparam DUL_8_TO_9   = 32'd3;    // 8->9: 3��
    localparam DUL_9_TO_10  = 32'd12;   // 9->10: 12��
    localparam DUL_10_TO_11 = 32'd9;    // 10->11: 9��
    localparam DUL_11_TO_12 = 32'd9;    // 11->12: 9��
    localparam DUL_12_TO_13 = 32'd15;   // 12->13: 15��
    localparam DUL_13_TO_14 = 32'd15;   // 13->14: 15��
    localparam DUL_14_FINAL = 32'd15;   // 14����: 15��
    
    // ��������ʱ��
    localparam BASE_DUL_LEN = 32'd10_000; // ��������ʱ��10ms
    localparam INIT_CNT = 16'd3000;    // ��ʼ���������
    
    // ���ͻ������ֵ
    localparam ERROR_THRESHOLD = 16'd100; // ���ͻ����ֵ���ӽ�2**15=32768��
    
    // �ڲ��ź�����
    reg                 pll_id;              // PLL�����ź�
    reg [PW-1:0]        r_phase_step;        // ��λ�����Ĵ���
    reg [4:0]           r_lg_coeff;          // ����ϵ���Ĵ���
    
    // �������״̬��
    reg [3:0]           r_stage;             // ������ƽ׶Σ�0-11��12���׶Σ�
    reg [15:0]          r_ice_cnt;           // ��ʼ������
    reg [31:0]          r_dul_cnt;           // ����ʱ�������
    reg [31:0]          r_current_dul_len;   // ��ǰ�׶γ���ʱ��
    reg [15:0]          r_prev_error_abs;    // ��һ����������ֵ
    
    
    
    // ���㵱ǰ������ֵ
    reg [15:0] current_error_abs;
    // �̶���λ����ֵ
    localparam FIXED_PHASE_STEP = 32'd429496;
    
    
    // ʵ����PLL����ģ��
    dblcordicpll #(
        .IW(IW),
        .PW(PW), 
        .OW(OW),
        .OPT_TRACK_FREQUENCY(1'b1),
        .OPT_FILTER(1'b1)
    ) u_pll_core (
        .i_clk        (clk),
        .i_reset      (~reset_n),        //�߸�λ
        .i_ld         (pll_id),     // Ӧ���ڸ�λ֮������
        .i_step       (r_phase_step),
        .i_ce         (enable_posedge), // ʹ��ad��������ΪPLLʹ��
        .i_input      (signal_in),   // ʹ��ͬ����������ź�
        .i_lgcoeff    (r_lg_coeff),
        .o_err        (phase_error),
        .o_phase      (output_phase),
        .pd_done      (pll_done) 
    );
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)begin
            pll_id <= 1;
        end else begin
            if (pll_id == 1) begin
                pll_id <= 0;
            end else if(r_error_jump)begin
               pll_id <= 1;
            end
        end
    end
    // ���ͻ�����߼�
    /*
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            r_prev_error_abs <= 16'd0;
            r_error_jump <= 1'b0;
        end else if (enable_posedge) begin  // ֻ��ad������ʱ���
            current_error_abs = phase_error;           
            // ������ͻ�䣺ֻ�����ս׶μ��
            if (r_stage == 4'd11 && (current_error_abs > phase_error + ERROR_THRESHOLD
                                     || current_error_abs < phase_error - ERROR_THRESHOLD)) begin
                r_error_jump <= 1'b0;
            end else begin
                r_error_jump <= 1'b0;
            end
            
            r_prev_error_abs <= current_error_abs;
        end
    end
    */
    // �������״̬�� - ������3��14��12���׶�
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            r_stage          <= 4'd0;
            r_ice_cnt        <= 16'd0;
            r_dul_cnt        <= 32'd0;
            r_lg_coeff       <= GAIN_3;
            r_current_dul_len <= BASE_DUL_LEN * DUL_3_TO_4;
        end else if (r_error_jump) begin
            // ���ͻ�䣺���õ���һ�׶�
            r_stage          <= 4'd0;
            r_ice_cnt        <= 16'd0;
            r_dul_cnt        <= 32'd0;
            r_lg_coeff       <= GAIN_3;
            r_current_dul_len <= BASE_DUL_LEN * DUL_3_TO_4;
        end else if (enable_posedge) begin  // ֻ��enable������ʱ����״̬��
            // ��ʼ�����׶�
            if (r_ice_cnt < INIT_CNT) begin
                r_ice_cnt <= r_ice_cnt + 16'd1;
                r_dul_cnt <= 32'd0;
            end else begin
                r_ice_cnt <= INIT_CNT + 16'd1; // ���̶ֹ�ֵ
                r_dul_cnt <= r_dul_cnt + 32'd1;
                
                // ״̬ת���߼� - ������3��14��12���׶�
                case (r_stage)
                    4'd0: begin // �׶�0������3
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd1;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_4;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_4_TO_5;
                        end
                    end
                    
                    4'd1: begin // �׶�1������4
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd2;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_5;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_5_TO_6;
                        end
                    end
                    
                    4'd2: begin // �׶�2������5
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd3;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_6;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_6_TO_7;
                        end
                    end
                    
                    4'd3: begin // �׶�3������6
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd4;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_7;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_7_TO_8;
                        end
                    end
                    
                    4'd4: begin // �׶�4������7
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd5;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_8;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_8_TO_9;
                        end
                    end
                    
                    4'd5: begin // �׶�5������8
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd6;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_9;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_9_TO_10;
                        end
                    end
                    
                    4'd6: begin // �׶�6������9
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd7;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_10;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_10_TO_11;
                        end
                    end
                    
                    4'd7: begin // �׶�7������10
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd8;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_11;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_11_TO_12;
                        end
                    end
                    
                    4'd8: begin // �׶�8������11
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd9;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_12;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_12_TO_13;
                        end
                    end
                    
                    4'd9: begin // �׶�9������12
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd10;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_13;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_13_TO_14;
                        end
                    end
                    
                    4'd10: begin // �׶�10������13
                        if (r_dul_cnt >= r_current_dul_len) begin
                            r_stage          <= 4'd11;
                            r_dul_cnt        <= 32'd0;
                            r_lg_coeff       <= GAIN_14;
                            r_current_dul_len <= BASE_DUL_LEN * DUL_14_FINAL;
                        end
                    end
                    
                    4'd11: begin // �׶�11������14�����ս׶Σ�
                        // ���ֵ�ǰ���棬�����л�
                        // �ȴ����ͻ��ǿ�Ƹ�λ
                    end
                    
                    default: begin
                        r_stage          <= 4'd0;
                        r_lg_coeff       <= GAIN_3;
                        r_current_dul_len <= BASE_DUL_LEN * DUL_3_TO_4;
                    end
                endcase
            end
        end
    end
    
    // ��λ�������ã��̶�ֵ��
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            r_phase_step <= FIXED_PHASE_STEP;
        end else begin
            r_phase_step <= FIXED_PHASE_STEP; // ���̶ֹ�
        end
    end

endmodule