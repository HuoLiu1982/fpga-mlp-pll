`timescale 1ns / 1ps

module lmlp_top (
    input  wire        clk_27M,
    input  wire        clk_135M,//�������135M,ʵ������ʹ��100M����pll����ʱ���Լ�adcʱ��ͳһ
    input  wire [15:0] ad_data_in,
    input  wire        rst_n,
    output reg [1:0]   mlp_prediction,
    output reg         mlp_done,
    output wire        uart_tx
);

/* -------------------------------------------------
 * 1MHz ����ʱ�� - �����汾
 * -------------------------------------------------*/
parameter DIVIDER = 100;
parameter CNT_MAX = DIVIDER/2 - 1;

reg clk_1M;
reg [7:0] clk_cnt;
reg clk_1M_prev;
reg pulse_ad;

always @(posedge clk_135M or negedge rst_n) begin
    if(!rst_n) begin
        clk_cnt <= 8'd0;
        clk_1M <= 1'b0;
        clk_1M_prev <= 1'b0;
        pulse_ad <= 1'b0;
    end else begin
        clk_1M_prev <= clk_1M;
        
        if(clk_cnt == CNT_MAX) begin
            clk_1M <= ~clk_1M;
            clk_cnt <= 8'd0;
        end else begin
            clk_cnt <= clk_cnt + 8'd1;
        end
        
        pulse_ad <= (clk_1M && !clk_1M_prev);
    end
end


/* -------------------------------------------------
 * �ϵ���ʱ��no��
 * -------------------------------------------------*/
reg        pwok;

always @(posedge clk_27M or negedge rst_n) begin
    if (!rst_n) begin
        pwok  <= 1;
    end
end

/* -------------------------------------------------
 * ADC�����͹�һ������
 * -------------------------------------------------*/
reg [10:0] addr;
reg        sample_done;
reg [15:0]  ad_buffer [0:63];
wire [15:0]  sample_data;
reg signed [31:0] normalized_data [0:63];

// Q10.22��ʽ����
localparam Q_FRAC_BITS = 22;
localparam Q_SCALE = 1 << Q_FRAC_BITS;

// ADC��һ��ϵ����1/255 in Q10.22 = 2^22 / 255���ĳ�1/2**16
localparam NORM_COEFF = 32'h00000040;

// ADC����״̬��
reg [1:0] adc_state;
localparam ADC_IDLE = 2'd0;
localparam ADC_SAMPLING = 2'd1;
localparam ADC_NORMALIZING = 2'd2;
localparam ADC_DONE = 2'd3;

reg [5:0] norm_addr;
reg [47:0] temp_product;  // 47λ�м���
reg signed [31:0] final_value;
integer i, j, k;
reg sample_en;
wire sam_done;
sample sample_uut(
    .clk_100M(clk_135M),
    .rst_n(rst_n),
    .enable(sample_en),
    .adc_dai_A(ad_data_in),
    .done(sam_done),
    .signal_tem(sample_data),//16λ
    .signal_out()//8λ
);

// ADC�����͹�һ������״̬��
always @(posedge clk_135M or negedge rst_n) begin
    if (!rst_n) begin
        adc_state <= ADC_IDLE;
        addr <= 0;
        norm_addr <= 0;
        sample_done <= 0;
        sample_en <= 0;
        // ��ʼ��������
        for (i = 0; i < 64; i = i + 1) begin
            ad_buffer[i] <= 0;
            normalized_data[i] <= 0;
        end
        $display("[ADC] ADC״̬����λ");
    end else if (pwok) begin  // ֻ���ϵ���ɺ������
        case(adc_state)
            ADC_IDLE: begin
                if (!sample_done) begin
                    adc_state <= ADC_SAMPLING;
                    sample_en <= 1;
                    addr <= 0;
                    $display("[ADC] ��ʼ����������ADC_SAMPLING״̬");
                end
            end
            
            ADC_SAMPLING: begin                        
                if (sam_done) begin
                    sample_en <= 0;
                    ad_buffer[addr] <= sample_data;
                    
                    if (addr == 63) begin
                        adc_state <= ADC_NORMALIZING;
                        addr <= 0;
                        norm_addr <= 0;
                    end else begin
                        addr <= addr + 1'd1;
                    end
                end
            end
            
            ADC_NORMALIZING: begin
                // �޷��ų˷�
                temp_product = ad_buffer[norm_addr] * NORM_COEFF;
                
                // ȷ���������ȷ�ķ�Χ�ڲ�ת��Ϊ�з���
                if (temp_product[47:32] != 16'b0) begin
                    // �����λ��Ϊ0��˵�������ʹ�����ֵ
                    final_value = 32'h3FFFFFF;  // �ӽ�1.0��Q10.22ֵ
                end else begin
                    // ���������ȡ��32λ��ȷ��������
                    final_value = {1'b0, temp_product[30:0]};  // ȷ������λΪ0
                end
                
                normalized_data[norm_addr] <= final_value;

                
                if (norm_addr == 63) begin
                    adc_state <= ADC_DONE;
                    sample_done <= 1;
                end else begin
                    norm_addr <= norm_addr + 1'd1;
                end
            end
            
            ADC_DONE: begin
                // �������״̬
            end
            
            default: begin
                adc_state <= ADC_IDLE;
                $display("[ADC] ���󣺽���δ֪״̬������IDLE");
            end
        endcase
    end else begin
        // �ϵ�δ��ɣ����ָ�λ״̬
        adc_state <= ADC_IDLE;
        sample_done <= 0;
    end
end
/* -------------------------------------------------
 * 5. MLP�������棨������ROM��ȡ�ͳ˷���
 * -------------------------------------------------*/
// �������ò���
localparam INPUT_SIZE = 64;
localparam HIDDEN_LAYER_1_SIZE = 32;
localparam HIDDEN_LAYER_2_SIZE = 16;
localparam OUTPUT_SIZE = 4;
// ����״̬��
reg [3:0] mlp_state;
reg [10:0] mlp_counter;
reg signed [63:0] mlp_mac_accumulator;  // ��Ϊ64λ��ֹ���
reg [4:0] mlp_neuron_idx;
reg [5:0] mlp_input_idx;

// �����ˮ�߿��ƼĴ���
reg pipeline_busy;

// �м���
reg signed [31:0] mlp_layer1_out [0:31];
reg signed [31:0] mlp_layer2_out [0:15];
reg signed [31:0] mlp_output_out [0:3];
reg [31:0] current_scale, current_shift;
reg signed [31:0] temp_relu;
reg signed [63:0] temp_mac;  // ��Ϊ64λ
reg signed [31:0] temp_bn;
reg signed [31:0] temp_bias;
// ������
reg [31:0] mlp_confidence;


// ״̬����
localparam MLP_IDLE = 4'd0;
localparam MLP_LAYER1_MAC = 4'd1;
localparam MLP_LAYER1_BIAS = 4'd2;
localparam MLP_LAYER1_BN = 4'd3;
localparam MLP_LAYER1_RELU = 4'd4;
localparam MLP_LAYER2_MAC = 4'd5;
localparam MLP_LAYER2_BIAS = 4'd6;
localparam MLP_LAYER2_BN = 4'd7;
localparam MLP_LAYER2_RELU = 4'd8;
localparam MLP_OUTPUT_MAC = 4'd9;
localparam MLP_OUTPUT_BIAS = 4'd10;
localparam MLP_FIND_MAX = 4'd11;
localparam MLP_DONE = 4'd12;

// ROM�ӿڣ�����layer1Ȩ�أ�
reg [10:0] rom_addr;
wire signed[31:0] rom_data;
rom_weights u_rom_weights (
  .addr(rom_addr),          // input [10:0]
  .clk(clk_135M),           // input
  .rst(!rst_n),             // input
  .rd_data(rom_data)        // output [31:0]
);

// LUT�ӿ�
wire signed[31:0] layer1_bias_data;
wire signed[31:0] layer2_weight_data;
wire signed[31:0] layer2_bias_data;
wire signed[31:0] output_weight_data;
wire signed[31:0] output_bias_data;
wire signed[31:0] bn1_scale_data;
wire signed[31:0] bn1_shift_data;
wire signed[31:0] bn2_scale_data;
wire signed[31:0] bn2_shift_data;

// ʵ����LUTģ��
layer1_bias_lut u_layer1_bias(.addr(mlp_neuron_idx), .data(layer1_bias_data));
layer2_weight_lut u_layer2_weight(.addr(rom_addr[9:0]), .data(layer2_weight_data));
layer2_bias_lut u_layer2_bias(.addr(mlp_neuron_idx), .data(layer2_bias_data));
output_weight_lut u_output_weight(.addr(rom_addr[5:0]), .data(output_weight_data));
output_bias_lut u_output_bias(.addr(mlp_neuron_idx), .data(output_bias_data));
bn1_scale_lut u_bn1_scale(.addr(mlp_neuron_idx), .data(bn1_scale_data));
bn1_shift_lut u_bn1_shift(.addr(mlp_neuron_idx), .data(bn1_shift_data));
bn2_scale_lut u_bn2_scale(.addr(mlp_neuron_idx), .data(bn2_scale_data));
bn2_shift_lut u_bn2_shift(.addr(mlp_neuron_idx), .data(bn2_shift_data));

// ROM��ȡ��ˮ�߿���
reg [1:0] rom_read_state;
reg signed [31:0] rom_data_reg;
reg signed [31:0] normalized_data_reg;
reg signed [31:0] layer1_out_reg;
reg        rom_read_valid;
reg signed [31:0] layer2_out_reg;
// �˷�����ˮ��
reg signed [63:0] multiply_result;
reg        multiply_valid;
reg [1:0]  multiply_state;

localparam ROM_READ_IDLE = 2'd0;
localparam ROM_READ_SETUP = 2'd1;
localparam ROM_READ_FETCH = 2'd2;

localparam MULTIPLY_IDLE = 2'd0;
localparam MULTIPLY_EXECUTE = 2'd1;

// ��������ź�
reg multiply_busy;           // �˷���æµ��־
reg [15:0] pending_rom_addr; // �������ROM��ַ


// ROM��ȡ״̬�� - ��ȫ��д
always @(posedge clk_135M or negedge rst_n) begin
    if (!rst_n) begin
        rom_read_state <= ROM_READ_IDLE;
        rom_read_valid <= 0;
        rom_data_reg <= 0;
        normalized_data_reg <= 0;
        layer1_out_reg <= 0;
        layer2_out_reg <= 0;
        multiply_busy <= 0;
        pending_rom_addr <= 0;
        $display("[ROM_READ] ROM��ȡ״̬����λ");
    end else begin
        rom_read_valid <= 0;
        
        case(rom_read_state)
            ROM_READ_IDLE: begin
                if ((mlp_state == MLP_LAYER1_MAC || mlp_state == MLP_LAYER2_MAC || 
                     mlp_state == MLP_OUTPUT_MAC) && !multiply_busy) begin
                    // ������ǰ��ַ�������ȡ
                    pending_rom_addr <= rom_addr;
                    rom_read_state <= ROM_READ_SETUP;
                    $display("[ROM_READ_IDLE] ����ROM��ȡ����ַ=%d��MLP״̬=%d", rom_addr, mlp_state);
                end
            end
            
            ROM_READ_SETUP: begin
                // ȷ��ROM��ַ�ȶ�
                if (rom_addr == pending_rom_addr) begin
                    // ׼����������
                    if (mlp_state == MLP_LAYER1_MAC) begin
                        normalized_data_reg <= normalized_data[mlp_input_idx];
                        $display("[ROM_READ_SETUP] L1_MAC: ��ַ=%d, ��һ������=%h", 
                                mlp_input_idx, normalized_data[mlp_input_idx]);
                    end else if (mlp_state == MLP_LAYER2_MAC) begin
                        layer1_out_reg <= mlp_layer1_out[mlp_input_idx];
                        $display("[ROM_READ_SETUP] L2_MAC: ��ַ=%d, ��1���=%h", 
                                mlp_input_idx, mlp_layer1_out[mlp_input_idx]);
                    end else if (mlp_state == MLP_OUTPUT_MAC) begin
                        layer2_out_reg <= mlp_layer2_out[mlp_input_idx];
                        $display("[ROM_READ_SETUP] OUT_MAC: ��ַ=%d, ��2���=%h", 
                                mlp_input_idx, mlp_layer2_out[mlp_input_idx]);
                    end
                    rom_read_state <= ROM_READ_FETCH;
                end else begin
                    // ��ַ�Ѹı䣬���¿�ʼ
                    $display("[ROM_READ_SETUP] ��ַ�ı䣬���¿�ʼ");
                    rom_read_state <= ROM_READ_IDLE;
                end
            end
            
            ROM_READ_FETCH: begin
                // ��ȡROM���ݲ����Ϊ��Ч
                rom_data_reg <= rom_data;
                rom_read_valid <= 1;
                multiply_busy <= 1; // ��ǳ˷�����ʼ����
                rom_read_state <= ROM_READ_IDLE;
                $display("[ROM_READ_FETCH] ��ȡROM����=%h����ַ=%d", rom_data, pending_rom_addr);
            end
        endcase
        
        // �˷����ʱ���æµ��־
        if (multiply_valid) begin
            multiply_busy <= 0;
            $display("[ROM_READ] �˷���ɣ����æµ��־");
        end
    end
end

// �˷���״̬��
always @(posedge clk_135M or negedge rst_n) begin
    if (!rst_n) begin
        multiply_result <= 0;
        multiply_valid <= 0;
        multiply_state <= MULTIPLY_IDLE;
        $display("[MULTIPLY] �˷�����ˮ�߸�λ");
    end else begin
        multiply_valid <= 0;
        
        case(multiply_state)
            MULTIPLY_IDLE: begin
                if (rom_read_valid && !multiply_valid) begin
                    multiply_state <= MULTIPLY_EXECUTE;
                    
                    // ִ�г˷�
                    if (mlp_state == MLP_LAYER1_MAC) begin
                        multiply_result <= rom_data_reg * normalized_data_reg;
                        $display("[MULTIPLY] L1_MAC: ROM����=%h * ��һ������=%h", 
                                rom_data_reg, normalized_data_reg);
                    end else if (mlp_state == MLP_LAYER2_MAC) begin
                        multiply_result <= layer2_weight_data * layer1_out_reg;
                        $display("[MULTIPLY] L2_MAC: Ȩ��=%h * ��1���=%h", 
                                layer2_weight_data, layer1_out_reg);
                    end else if (mlp_state == MLP_OUTPUT_MAC) begin
                        multiply_result <= output_weight_data * layer2_out_reg;
                        $display("[MULTIPLY] OUT_MAC: Ȩ��=%h * ��2���=%h", 
                                output_weight_data, layer2_out_reg);
                    end
                end
            end
            
            MULTIPLY_EXECUTE: begin
                multiply_valid <= 1;
                multiply_state <= MULTIPLY_IDLE;
                $display("[MULTIPLY] �˷���ɣ����=%h", multiply_result);
            end
        endcase
    end
end


// ��ȡQ10.22���
function signed [31:0] extract_q10_22;
    input signed [63:0] product;
    reg signed [31:0] result;
    begin
        // ���ƫ������������
        product = product + (1 << (Q_FRAC_BITS - 1));
        result = product >>> Q_FRAC_BITS;  // ����22λ�õ�Q10.22
        $display("[EXTRACT_Q10_22] ����˻�=%h, ������=%h", product, result);
        extract_q10_22 = result;
    end
endfunction

// 64λ��32λ���з��ű��ʹ���
function signed [31:0] saturate_64_to_32;
    input signed [63:0] value;
    begin
        if (value > $signed(64'sh000000007FFFFFFF)) begin
            // ����32λ�з������ֵ�����͵����ֵ
            saturate_64_to_32 = 32'sh7FFFFFFF;
            $display("[SATURATE] 64λֵ=%h ����32λ�����ֵ�����͵�7FFFFFFF", value);
        end else if (value < $signed(64'shFFFFFFFF80000000)) begin
            // С��32λ�з�����Сֵ�����͵���Сֵ
            saturate_64_to_32 = 32'sh80000000;
            $display("[SATURATE] 64λֵ=%h ����32λ����Сֵ�����͵�80000000", value);
        end else begin
            // ��32λ��Χ�ڣ�ֱ�ӽض�
            saturate_64_to_32 = value[31:0];
            $display("[SATURATE] 64λֵ=%h ��32λ��Χ�ڣ��ض�Ϊ=%h", value, value[31:0]);
        end
    end
endfunction

// ������ReLU�����
function signed [31:0] relu_fixed;
    input signed [31:0] x;
    begin
        if (x < 0) begin
            $display("[RELU] ����=%h (����), ���=0", x);
            relu_fixed = 0;
        end else begin
            $display("[RELU] ����=%h (����), ������ֲ���", x);
            relu_fixed = x;
        end      
    end
endfunction

// �Ľ���BatchNormʵ��
function signed [31:0] batchnorm_simple;
    input signed [31:0] x;
    input signed [31:0] scale;
    input signed [31:0] shift;
    reg signed [63:0] scaled;
    reg signed [63:0] rounded;
    begin
        scaled = $signed(x) * $signed(scale);
        // ���õ����봦��
        rounded = scaled + (1 << (Q_FRAC_BITS - 1));
        batchnorm_simple = (rounded >>> Q_FRAC_BITS) + shift;
        
        $display("[IMPROVED_BN] x=%h, scale=%h, scaled=%h, result=%h", 
                 x, scale, scaled, batchnorm_simple);
    end
endfunction

// ��ʱ����ͬ�������sample_done�������أ�3MHz -> 135MHz��
reg sample_done_sync1, sample_done_sync2, sample_done_sync3;
wire sample_done_rising;

always @(posedge clk_135M or negedge rst_n) begin
    if (!rst_n) begin
        sample_done_sync1 <= 0;
        sample_done_sync2 <= 0;
        sample_done_sync3 <= 0;
    end else begin
        sample_done_sync1 <= sample_done;
        sample_done_sync2 <= sample_done_sync1;
        sample_done_sync3 <= sample_done_sync2;
    end
end
assign sample_done_rising = sample_done_sync2 && !sample_done_sync3;

// MLP����״̬����135MHzʱ�ӣ�
always @(posedge clk_135M or negedge rst_n) begin
    if (!rst_n) begin
        mlp_state <= MLP_IDLE;
        mlp_counter <= 0;
        mlp_done <= 0;
        mlp_prediction <= 0;
        mlp_confidence <= 0;
        rom_addr <= 0;
        mlp_mac_accumulator <= 0;
        mlp_neuron_idx <= 0;
        mlp_input_idx <= 0;
        pipeline_busy <= 0;
        // ��ʼ������
        for (i = 0; i < 32; i = i + 1) mlp_layer1_out[i] <= 0;
        for (j = 0; j < 16; j = j + 1) mlp_layer2_out[j] <= 0;
        for (k = 0; k < 4; k = k + 1) mlp_output_out[k] <= 0;
        
        $display("[MLP] MLP״̬����λ");
    end else begin
        case(mlp_state)
            MLP_IDLE: begin
                if (sample_done_rising) begin
                    mlp_state <= MLP_LAYER1_MAC;
                    mlp_counter <= 0;
                    mlp_neuron_idx <= 0;
                    mlp_input_idx <= 0;
                    rom_addr <= 0;
                    mlp_mac_accumulator <= 0;
                    $display("[MLP] ��ʼ��������MLP_LAYER1_MAC״̬");
                end
                mlp_done <= 0;
            end
            
            MLP_LAYER1_MAC: begin
                // ��ǰ����ROM��ַ��ȷ����ROM��ȡ��ʼǰ��ַ���ȶ�
                if (!pipeline_busy && rom_read_state == ROM_READ_IDLE) begin
                    rom_addr <= (mlp_neuron_idx * INPUT_SIZE) + mlp_input_idx;
                    pipeline_busy <= 1;  // �����ˮ��æµ
                    $display("[MLP_LAYER1_MAC] ����ROM��ַ=%d", (mlp_neuron_idx * INPUT_SIZE) + mlp_input_idx);
                end
                if (mlp_counter < 2048) begin                   
                    if (multiply_valid) begin
                        // �ۼӳ˷���� - ʹ��64λ�ۼ���
                        temp_mac = mlp_mac_accumulator + $signed(extract_q10_22(multiply_result));
                        //temp_mac = mlp_mac_accumulator + $signed(multiply_result);
                        mlp_mac_accumulator <= temp_mac;
                        
                        $display("[MLP_LAYER1_MAC] MAC����: ������=%d, ��Ԫ=%d, ����=%d, ���ۼ���=%h, ���ۼ���=%h", 
                                 mlp_counter, mlp_neuron_idx,mlp_input_idx, mlp_mac_accumulator, temp_mac);
                        
                        mlp_input_idx <= mlp_input_idx + 1;
                        pipeline_busy <= 0;  // ���æµ��־������������һ�ζ�ȡ
                        if (mlp_input_idx == 63) begin
                            // ��ɵ�ǰ��Ԫ��ȫ������
                            mlp_state <= MLP_LAYER1_BIAS;
                            mlp_input_idx <= 0;
                            $display("[MLP] ��1 MAC��ɣ�����BIAS״̬");
                        end else begin
                            // ׼����һ������
                            mlp_counter <= mlp_counter + 1;
                            $display("[MLP_LAYER1_MAC] ׼����һ�����룬�¼�����=%d", mlp_counter + 1);
                        end
                    end
                 end else begin
                        // ��ֹ����
                        mlp_state <= MLP_LAYER1_BIAS;
                        mlp_input_idx <= 0;
                        pipeline_busy <= 0;  // ���æµ��־
                        $display("[MLP] ���棺���������ޣ�ǿ�ƽ���BIAS״̬");
                end
            end
            MLP_LAYER1_BIAS: begin
                // ���ƫ�� - ʹ�ñ��ʹ���64λת��Ϊ32λ
                rom_addr <= mlp_neuron_idx;
                
                // ��ƫ�÷�����չΪ64λ��Ȼ�����ۼ�����ӣ������б��ʹ���
                temp_mac = mlp_mac_accumulator + {{32{layer1_bias_data[31]}}, layer1_bias_data};
                temp_bias = saturate_64_to_32(temp_mac);
                mlp_layer1_out[mlp_neuron_idx] <= temp_bias;
                mlp_mac_accumulator <= 0;
                
                $display("[MLP_LAYER1_BIAS] ��Ԫ=%d, MAC���=%h, ƫ��=%h, �������=%h", 
                         mlp_neuron_idx, mlp_mac_accumulator, layer1_bias_data, mlp_layer1_out[mlp_neuron_idx]);
                
                // ������һ����Ԫ����ʼ��ַ
                mlp_counter <= (mlp_neuron_idx + 1) * 64;
                mlp_input_idx <= 0;
                pipeline_busy <= 0;
                mlp_mac_accumulator <= 0;
                if (mlp_neuron_idx == 31) begin
                    // ������Ԫ�������
                    mlp_state <= MLP_LAYER1_BN;
                            mlp_neuron_idx <= 0;
                            mlp_input_idx <= 0;
                            pipeline_busy <= 0;  // ���æµ��־
                    rom_addr <= 0;
                    $display("[MLP] ��1ƫ����ɣ�����BN״̬");
                end else begin
                    // ������һ����Ԫ
                    mlp_neuron_idx <= mlp_neuron_idx + 1;
                    mlp_state <= MLP_LAYER1_MAC;
                    $display("[MLP] ������һ����Ԫ: %d", mlp_neuron_idx + 1);
                end
            end
            
            MLP_LAYER1_BN: begin
                // ����BN������ַ
                rom_addr <= mlp_neuron_idx;
                
                // ʹ�üĴ����ݴ�BN��������������߼��ӳ�               
                current_scale = bn1_scale_data;
                current_shift = bn1_shift_data;
                
                $display("[MLP_LAYER1_BN] ��Ԫ=%d, ����=%h, scale=%h, shift=%h", 
                         mlp_neuron_idx, mlp_layer1_out[mlp_neuron_idx], current_scale, current_shift);
                
                temp_bn = batchnorm_simple(
                    mlp_layer1_out[mlp_neuron_idx],
                    current_scale,
                    current_shift
                );
                mlp_layer1_out[mlp_neuron_idx] <= temp_bn;
                $display("[MLP_LAYER1_BN] BN�����=%h", temp_bn);
                
                mlp_neuron_idx <= mlp_neuron_idx + 1;
                
                if (mlp_neuron_idx == 31) begin
                    mlp_state <= MLP_LAYER1_RELU;
                    mlp_neuron_idx <= 0;
                    rom_addr <= 0;
                    $display("[MLP] ��1 BN��ɣ�����RELU״̬");
                end
            end
            
            MLP_LAYER1_RELU: begin
                // ReLU����һ���������������Ԫ
                for (i = 0; i < 32; i = i + 1) begin
                    temp_relu = relu_fixed(mlp_layer1_out[i]);
                    mlp_layer1_out[i] <= temp_relu;
                    $display("[MLP_LAYER1_RELU] ��Ԫ=%d, ReLU��=%h", i, temp_relu);
                end
                mlp_state <= MLP_LAYER2_MAC;
                mlp_neuron_idx <= 0;
                mlp_input_idx <= 0;
                mlp_counter <= 0;
                rom_addr <= 0;
                $display("[MLP] ��1 RELU��ɣ������2 MAC״̬");
            end
            
            MLP_LAYER2_MAC: begin
                if (mlp_counter < 512) begin
                    if (!pipeline_busy && rom_read_state == ROM_READ_IDLE) begin
                        rom_addr <= mlp_counter;
                        pipeline_busy <= 1;
                        $display("[MLP_LAYER2_MAC] ����ROM��ȡ����ַ=%d", mlp_counter);
                    end
                    
                    if (multiply_valid) begin
                        // �ۼӳ˷���� - ʹ��64λ�ۼ���
                        temp_mac = mlp_mac_accumulator + $signed(extract_q10_22(multiply_result));
                        //temp_mac = mlp_mac_accumulator + $signed(multiply_result);
                        mlp_mac_accumulator <= temp_mac;
                        
                        $display("[MLP_LAYER2_MAC] MAC����: ������=%d, ��Ԫ=%d,����=%d, ���ۼ���=%h, ���ۼ���=%h", 
                                 mlp_counter, mlp_neuron_idx,mlp_input_idx, mlp_mac_accumulator, temp_mac);
                        
                        mlp_input_idx <= mlp_input_idx + 1;
                        
                        if (mlp_input_idx == 31) begin
                            mlp_state <= MLP_LAYER2_BIAS;
                            mlp_input_idx <= 0;
                            pipeline_busy <= 0;  // ���æµ��־
                            $display("[MLP] ��2 MAC��ɣ�����BIAS״̬");
                        end else begin
                            mlp_counter <= mlp_counter + 1;
                            pipeline_busy <= 0;
                            $display("[MLP_LAYER2_MAC] ׼����һ�����룬�¼�����=%d", mlp_counter + 1);
                        end
                    end
                end else begin
                    mlp_state <= MLP_LAYER2_BIAS;
                            mlp_input_idx <= 0;
                            pipeline_busy <= 0;  // ���æµ��־
                    $display("[MLP] ���棺���������ޣ�ǿ�ƽ���BIAS״̬");
                end
            end           
            MLP_LAYER2_BIAS: begin
                rom_addr <= mlp_neuron_idx;
                // ��ƫ�÷�����չΪ64λ��Ȼ�����ۼ�����ӣ������б��ʹ���
                temp_mac = mlp_mac_accumulator + {{32{layer2_bias_data[31]}}, layer2_bias_data};
                temp_bias = saturate_64_to_32(temp_mac);
                mlp_layer2_out[mlp_neuron_idx] <= temp_bias;
                mlp_mac_accumulator <= 0;
                
                $display("[MLP_LAYER2_BIAS] ��Ԫ=%d, MAC���=%h, ƫ��=%h, �������=%h", 
                         mlp_neuron_idx, mlp_mac_accumulator, layer2_bias_data, mlp_layer2_out[mlp_neuron_idx]);
                
                // ������һ����Ԫ����ʼ��ַ
                mlp_counter <= (mlp_neuron_idx + 1) * 32;
                mlp_input_idx <= 0;
                pipeline_busy <= 0;
                mlp_mac_accumulator <= 0;
                if (mlp_neuron_idx == 15) begin
                    mlp_state <= MLP_LAYER2_BN;
                    mlp_neuron_idx <= 0;
                    rom_addr <= 0;
                    $display("[MLP] ��2ƫ����ɣ�����BN״̬");
                end else begin
                    mlp_neuron_idx <= mlp_neuron_idx + 1;
                    mlp_state <= MLP_LAYER2_MAC;
                    $display("[MLP] ������һ����Ԫ: %d", mlp_neuron_idx + 1);
                end
            end
            
            MLP_LAYER2_BN: begin
                // ������ַ����
                rom_addr <= mlp_neuron_idx[3:0];  // ֱ��ʹ��4λ��ַ
                current_scale = bn2_scale_data;
                current_shift = bn2_shift_data;
                
                $display("[MLP_LAYER2_BN] ��Ԫ=%d, ����=%h, scale=%h, shift=%h", 
                         mlp_neuron_idx, mlp_layer2_out[mlp_neuron_idx], current_scale, current_shift);
                
                temp_bn = batchnorm_simple(
                    mlp_layer2_out[mlp_neuron_idx],
                    current_scale,
                    current_shift
                );
                mlp_layer2_out[mlp_neuron_idx] <= temp_bn;
                $display("[MLP_LAYER2_BN] BN�����=%h", temp_bn);
                
                mlp_neuron_idx <= mlp_neuron_idx + 1;
                
                if (mlp_neuron_idx == 15) begin
                    mlp_state <= MLP_LAYER2_RELU;
                    mlp_neuron_idx <= 0;
                    rom_addr <= 0;
                    $display("[MLP] ��2 BN��ɣ�����RELU״̬");
                end
            end
            
            MLP_LAYER2_RELU: begin
                // ReLU����һ���������������Ԫ
                for (i = 0; i < 16; i = i + 1) begin
                    temp_relu = relu_fixed(mlp_layer2_out[i]);
                    mlp_layer2_out[i] <= temp_relu;
                    $display("[MLP_LAYER2_RELU] ��Ԫ=%d, ReLU��=%h", i, temp_relu);
                end
                mlp_state <= MLP_OUTPUT_MAC;
                mlp_neuron_idx <= 0;
                mlp_input_idx <= 0;
                mlp_counter <= 0;
                rom_addr <= 0;
                $display("[MLP] ��2 RELU��ɣ����������MAC״̬");
            end
            
            MLP_OUTPUT_MAC: begin
                if (mlp_counter < 64) begin
                    if (rom_read_state == ROM_READ_IDLE) begin
                        rom_addr <= mlp_counter;
                    end
                    
                    if (multiply_valid) begin
                        // �ۼӳ˷���� - ʹ��64λ�ۼ���
                        temp_mac = mlp_mac_accumulator + $signed(extract_q10_22(multiply_result));
                        //temp_mac = mlp_mac_accumulator + $signed(multiply_result);
                        mlp_mac_accumulator <= temp_mac;
                        mlp_input_idx <= mlp_input_idx + 1;
                        mlp_counter <= mlp_counter + 1;
                        
                        $display("[MLP_OUTPUT_MAC] MAC����: ������=%d, ��Ԫ=%d,�ۼ���=%h,���ۼ���=%h",
                            mlp_counter, mlp_neuron_idx, mlp_mac_accumulator,temp_mac);
                        
                        if (mlp_input_idx == 15) begin
                            mlp_state <= MLP_OUTPUT_BIAS;
                            mlp_input_idx <= 0;
                            $display("[MLP] ����� MAC��ɣ�����BIAS״̬");
                        end else begin
                            rom_addr <= mlp_counter + 1;
                        end
                    end
                end else begin
                    // ��ֹ����
                    mlp_state <= MLP_OUTPUT_BIAS;
                    $display("[MLP] ���棺���������ޣ�ǿ�ƽ���BIAS״̬");
                end
            end
            
            MLP_OUTPUT_BIAS: begin
                // ��ƫ�÷�����չΪ64λ��Ȼ�����ۼ�����ӣ������б��ʹ���
                temp_mac = mlp_mac_accumulator + {{32{output_bias_data[31]}}, output_bias_data};
                temp_bias = saturate_64_to_32(temp_mac);
                mlp_output_out[mlp_neuron_idx] <= temp_bias;
                mlp_mac_accumulator <= 0;
                
                $display("[MLP_OUTPUT_BIAS] �����Ԫ=%d, MAC���=%h, ƫ��=%h, �������=%h", 
                         mlp_neuron_idx, mlp_mac_accumulator, output_bias_data, mlp_output_out[mlp_neuron_idx]);
                
                mlp_neuron_idx <= mlp_neuron_idx + 1;
                
                if (mlp_neuron_idx == 3) begin
                    mlp_state <= MLP_FIND_MAX;
                    mlp_neuron_idx <= 0;
                    $display("[MLP] �����ƫ����ɣ�����FIND_MAX״̬");
                end else begin
                    mlp_state <= MLP_OUTPUT_MAC;
                    mlp_counter <= (mlp_neuron_idx + 1) * 16;
                    mlp_input_idx <= 0;
                    $display("[MLP] ������һ�������Ԫ: %d", mlp_neuron_idx + 1);
                end
            end
            
            MLP_FIND_MAX: begin
                // �ҵ����ֵ��ΪԤ����
                $display("[MLP_FIND_MAX] ���ֵ: [0]=%h, [1]=%h, [2]=%h, [3]=%h", 
                         mlp_output_out[0], mlp_output_out[1], mlp_output_out[2], mlp_output_out[3]);
                
                if (mlp_output_out[0] >= mlp_output_out[1] && 
                    mlp_output_out[0] >= mlp_output_out[2] && 
                    mlp_output_out[0] >= mlp_output_out[3]) begin
                    mlp_prediction <= 2'b00; // ���Ҳ�
                    mlp_confidence <= mlp_output_out[0];
                    $display("[MLP_FIND_MAX] Ԥ����: ���Ҳ�, ���Ŷ�=%h", mlp_output_out[0]);
                end else if (mlp_output_out[1] >= mlp_output_out[0] && 
                           mlp_output_out[1] >= mlp_output_out[2] && 
                           mlp_output_out[1] >= mlp_output_out[3]) begin
                    mlp_prediction <= 2'b01; // ����
                    mlp_confidence <= mlp_output_out[1];
                    $display("[MLP_FIND_MAX] Ԥ����: ����, ���Ŷ�=%h", mlp_output_out[1]);
                end else if (mlp_output_out[2] >= mlp_output_out[0] && 
                           mlp_output_out[2] >= mlp_output_out[1] && 
                           mlp_output_out[2] >= mlp_output_out[3]) begin
                    mlp_prediction <= 2'b10; // ���ǲ�
                    mlp_confidence <= mlp_output_out[2];
                    $display("[MLP_FIND_MAX] Ԥ����: ���ǲ�, ���Ŷ�=%h", mlp_output_out[2]);
                end else begin
                    mlp_prediction <= 2'b11; // ����
                    mlp_confidence <= mlp_output_out[3];
                    $display("[MLP_FIND_MAX] Ԥ����: ����, ���Ŷ�=%h", mlp_output_out[3]);
                end
                mlp_state <= MLP_DONE;
            end
            
            MLP_DONE: begin
                mlp_done <= 1;
                $display("[MLP_DONE] MLP�������! Ԥ��=%b, ���Ŷ�=%h", mlp_prediction, mlp_confidence);
                // ����״ֱ̬���µĲ�����ʼ
                if (!sample_done_sync2) begin
                    mlp_state <= MLP_IDLE;
                    mlp_done <= 0;
                    $display("[MLP] ����IDLE״̬���ȴ���һ������");
                end
            end
            
            default: begin
                mlp_state <= MLP_IDLE;
                $display("[MLP] ���󣺽���δ֪״̬������IDLE");
            end
        endcase
    end
end
/* -------------------------------------------------
 * 6. UART���Ϳ��� - ��չ֧��MLP�����ӡ
 * -------------------------------------------------*/
reg [10:0] uart_cnt;
reg [7:0]  uart_data;
reg        uart_start_send;
reg        uart_sending;
reg        mlp_done_reg;
reg [2:0]  uart_state;
wire       mlp_done_rising;
// UART����״̬��
localparam UART_IDLE = 3'd0;
localparam UART_SEND_ADC_HEADER = 3'd1;
localparam UART_SEND_ADC_DATA = 3'd2;
localparam UART_SEND_MLP_HEADER = 3'd3;
localparam UART_SEND_MLP_RESULT = 3'd4;
localparam UART_SEND_CONFIDENCE = 3'd5;
localparam UART_DONE = 3'd6;
// ��ʱ����ͬ�������mlp_done�������أ�135MHz -> 27MHz��
// MLP�źſ�ʱ����ͬ����27MHz
reg mlp_done_sync_27M;
reg mlp_done_sync_27M_delay;
reg [1:0] mlp_prediction_sync_27M;
reg [31:0] mlp_confidence_sync_27M;

// ͬ��mlp_done�źŲ����������
always @(posedge clk_27M or negedge rst_n) begin
    if (!rst_n) begin
        mlp_done_sync_27M <= 0;
        mlp_done_sync_27M_delay <= 0;
        mlp_prediction_sync_27M <= 0;
        mlp_confidence_sync_27M <= 0;
    end else begin
        // ��һ��ͬ��
        mlp_done_sync_27M <= mlp_done;
        mlp_prediction_sync_27M <= mlp_prediction;
        mlp_confidence_sync_27M <= mlp_confidence;
        
        // �ڶ���ͬ�����ӳ����ڱ��ؼ��
        mlp_done_sync_27M_delay <= mlp_done_sync_27M;
    end
end

// ���ͬ�����mlp_done������
wire mlp_done_rising_sync = mlp_done_sync_27M && !mlp_done_sync_27M_delay;

// ����ֵת��Ϊʮ������ASCII�ַ�
function [7:0] byte_to_hex_ascii;
    input [7:0] data;
    input integer nibble; // 0: ��4λ, 1: ��4λ
    reg [3:0] nibble_data;
    begin
        nibble_data = (nibble == 0) ? data[7:4] : data[3:0];
        if (nibble_data <= 9)
            byte_to_hex_ascii = 8'h30 + nibble_data; // '0'-'9'
        else
            byte_to_hex_ascii = 8'h41 + (nibble_data - 10); // 'A'-'F'
    end
endfunction

// ��16λ��ֵת��Ϊʮ������ASCII�ַ�
function [7:0] word_to_hex_ascii;
    input [15:0] data;
    input integer nibble; // 0: ���4λ, 1: �θ�4λ, 2: �ε�4λ, 3: ���4λ
    reg [3:0] nibble_data;
    begin
        case(nibble)
            0: nibble_data = data[15:12];
            1: nibble_data = data[11:8];
            2: nibble_data = data[7:4];
            3: nibble_data = data[3:0];
            default: nibble_data = 4'b0;
        endcase
        if (nibble_data <= 9)
            word_to_hex_ascii = 8'h30 + nibble_data; // '0'-'9'
        else
            word_to_hex_ascii = 8'h41 + (nibble_data - 10); // 'A'-'F'
    end
endfunction

// �����Ŷ�ת��ΪASCII�ַ���
function [7:0] confidence_to_ascii;
    input [31:0] conf_q10_22;
    integer conf_int;
    begin
        // ��Q10.22ת��Ϊ0-100�������ٷֱ�
        conf_int = (conf_q10_22 * 100) >>> Q_FRAC_BITS;
        if (conf_int > 99) conf_int = 99;
        if (conf_int < 0) conf_int = 0;
        
        // ת��Ϊ��λASCII����
        if (conf_int >= 10) begin
            confidence_to_ascii = 8'h30 + (conf_int / 10);  // ʮλ
        end else begin
            confidence_to_ascii = 8'h30;  // ʮλΪ0
        end
    end
endfunction

// ��ȡ�����ַ���
function [7:0] get_type_char;
    input [1:0] pred;
    input integer pos;
    begin
        case(pred)
            2'b00: get_type_char = (pos == 0) ? "S" : (pos == 1) ? "I" : (pos == 2) ? "N" : " ";  // "SIN"
            2'b01: get_type_char = (pos == 0) ? "S" : (pos == 1) ? "Q" : (pos == 2) ? "U" : " ";  // "SQU"
            2'b10: get_type_char = (pos == 0) ? "T" : (pos == 1) ? "R" : (pos == 2) ? "I" : " ";  // "TRI"
            2'b11: get_type_char = (pos == 0) ? "O" : (pos == 1) ? "T" : (pos == 2) ? "H" : " ";  // "OTH"
            default: get_type_char = " ";
        endcase
    end
endfunction
integer conf_int;
// UART����״̬�� - �ϲ���ĵ���always��
always @(posedge clk_27M or negedge rst_n) begin
    if (!rst_n) begin
        uart_state <= UART_IDLE;
        uart_cnt <= 0;
        uart_data <= 0;
        uart_start_send <= 0;
        uart_sending <= 0;
    end else begin
        uart_start_send <= 0;
        
        // ����ѡ���߼� - ���ݵ�ǰ״̬�ͼ�����ѡ��Ҫ���͵�����
        case(uart_state)
            UART_SEND_ADC_HEADER: begin
                case(uart_cnt)
                    0: uart_data <= "A";
                    1: uart_data <= "D";
                    2: uart_data <= "C";
                    3: uart_data <= ":";
                    default: uart_data <= 0;
                endcase
            end
            
            UART_SEND_ADC_DATA: begin
                // ÿ��16λ���ݷ���4��ʮ�������ַ�
                case(uart_cnt[1:0])
                    0: uart_data <= word_to_hex_ascii(ad_buffer[uart_cnt[9:2]], 0); // ���4λ
                    1: uart_data <= word_to_hex_ascii(ad_buffer[uart_cnt[9:2]], 1); // �θ�4λ
                    2: uart_data <= word_to_hex_ascii(ad_buffer[uart_cnt[9:2]], 2); // �ε�4λ
                    3: uart_data <= word_to_hex_ascii(ad_buffer[uart_cnt[9:2]], 3); // ���4λ
                    default: uart_data <= 0;
                endcase
            end
            
            UART_SEND_MLP_HEADER: begin
                case(uart_cnt)
                    0: uart_data <= " ";
                    1: uart_data <= "M";
                    2: uart_data <= "L";
                    3: uart_data <= "P";
                    4: uart_data <= ":";
                    default: uart_data <= 0;
                endcase
            end
            
            UART_SEND_MLP_RESULT: begin
                uart_data <= get_type_char(mlp_prediction_sync_27M, uart_cnt);
            end
            
            UART_SEND_CONFIDENCE: begin
                case(uart_cnt)
                    0: uart_data <= " ";
                    1: uart_data <= confidence_to_ascii(mlp_confidence_sync_27M);  // ʮλ
                    2: begin
                        
                        conf_int = (mlp_confidence_sync_27M * 100) >>> Q_FRAC_BITS;
                        if (conf_int > 99) conf_int = 99;
                        if (conf_int < 0) conf_int = 0;
                        uart_data <= 8'h30 + (conf_int % 10);  // ��λ
                    end
                    3: uart_data <= "%";  // �ٷֱȷ���
                    4: uart_data <= "\r"; // �س�
                    5: uart_data <= "\n"; // ����
                    default: uart_data <= 0;
                endcase
            end
            
            default: uart_data <= 0;
        endcase
        
        // ״̬ת�ƿ����߼�
        if (uart_sending && uart_start_send) begin
            uart_start_send <= 0;  // ��������ź�
        end
        else if (uart_sending && tx_busy_falling) begin
            // ��ǰ�ַ�������ɣ�׼��������һ��
            case(uart_state)
                UART_SEND_ADC_HEADER: begin
                    if (uart_cnt < 3) begin
                        uart_cnt <= uart_cnt + 1;
                        uart_start_send <= 1;
                    end else begin
                        uart_state <= UART_SEND_ADC_DATA;
                        uart_cnt <= 0;
                        uart_start_send <= 1;  // ������ʼ����ADC����
                    end
                end
                
                UART_SEND_ADC_DATA: begin
                    if (uart_cnt < 255) begin  // 64��16λ���� �� 4�ַ� = 256
                        uart_cnt <= uart_cnt + 1;
                        uart_start_send <= 1;
                    end else begin
                        uart_state <= UART_SEND_MLP_HEADER;
                        uart_cnt <= 0;
                        uart_start_send <= 1;  // ������ʼ����MLPͷ��
                    end
                end
                
                UART_SEND_MLP_HEADER: begin
                    if (uart_cnt < 4) begin
                        uart_cnt <= uart_cnt + 1;
                        uart_start_send <= 1;
                    end else begin
                        uart_state <= UART_SEND_MLP_RESULT;
                        uart_cnt <= 0;
                        uart_start_send <= 1;  // ������ʼ����MLP���
                    end
                end
                
                UART_SEND_MLP_RESULT: begin
                    if (uart_cnt < 2) begin  // ����3���ַ���0,1,2
                        uart_cnt <= uart_cnt + 1;
                        uart_start_send <= 1;
                    end else begin
                        uart_state <= UART_SEND_CONFIDENCE;
                        uart_cnt <= 0;
                        uart_start_send <= 1;  // ������ʼ�������Ŷ�
                    end
                end
                
                UART_SEND_CONFIDENCE: begin
                    if (uart_cnt < 5) begin  // ����6���ַ���0-5
                        uart_cnt <= uart_cnt + 1;
                        uart_start_send <= 1;
                    end else begin
                        uart_state <= UART_DONE;
                        uart_sending <= 0;  // �������
                    end
                end
                
                default: begin
                    uart_state <= UART_IDLE;
                    uart_sending <= 0;
                end
            endcase
        end
        else if (!uart_sending && mlp_done_rising_sync) begin
            // ʹ��ͬ�����MLP����ź�����UART����
            uart_state <= UART_SEND_ADC_HEADER;
            uart_sending <= 1;
            uart_cnt <= 0;
            uart_start_send <= 1;  // ������ʼ����
            
            // ���õ�һ��Ҫ���͵�����
            uart_data <= "A";
        end
    end
end
// ���tx_busy�½���
reg tx_busy_reg;
always @(posedge clk_27M or negedge rst_n) begin
    if (!rst_n) begin
        tx_busy_reg <= 0;
    end else begin
        tx_busy_reg <= tx_busy;
    end
end
wire tx_busy_falling = (!tx_busy) && tx_busy_reg;

// UART����ģ��ʵ����
wire tx_busy;
uart_tx_only my_uart_tx (
    .clk        (clk_27M),
    .temp_data  (uart_data),
    .start_send (uart_start_send),
    .uart_tx    (uart_tx),
    .tx_busy    (tx_busy)
);
endmodule