module triangle_wave(
    input clk,
    input [31:0] phase,
    output reg signed [15:0] triangle_out
);

    // ֱ��ʹ����λ�ĸ�16λ��Ϊ����ӳ��
    wire [15:0] linear;
    assign linear = phase[31:16];
    
    // ���ǲ����ɣ��������λ����б��
    always @(posedge clk) begin
        if (phase[31] == 1'b0) begin
            // ǰ�����ڣ�����
            triangle_out <= {1'b0, linear[14:0]} - 16'd16384; // -16384 to +16383
        end else begin
            // ������ڣ��½�  
            triangle_out <= 16'd16384 - {1'b0, linear[14:0]}; // +16383 to -16384
        end
    end

endmodule