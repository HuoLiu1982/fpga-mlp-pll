module key_ctrl(
    input  wire clk,
    input  wire rst_n,
    input  wire key_in,        // �������루�͵�ƽ��Ч��
    output reg  key_short,     // �̰����������������壩
    output reg  key_long       // �������������������壩
   );

    parameter CLK_FREQ = 27_000_000;
    parameter DEBOUNCE_MS = 20;
    parameter HOLD_MS = 1000;

    parameter CNT_20MS = (CLK_FREQ/1000)*DEBOUNCE_MS;   // 20msȥ��
    parameter CNT_1S   = (CLK_FREQ/1000)*HOLD_MS;       // 1�볤���ж�

    reg key_sync0, key_sync1;
    reg key_state;          // ��ǰ�ȶ�����״̬
    reg [31:0] cnt_debounce;
    reg [31:0] cnt_hold;

    // ===================== �ź�ͬ����������̬�� =====================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            key_sync0 <= 1'b1;
            key_sync1 <= 1'b1;
        end else begin
            key_sync0 <= key_in;
            key_sync1 <= key_sync0;
        end
    end

    // ===================== 20msȥ���� =====================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cnt_debounce <= 0;
            key_state <= 1'b1; // ��ʼδ����
        end else begin
            if (key_sync1 != key_state) begin
                cnt_debounce <= cnt_debounce + 1;
                if (cnt_debounce >= CNT_20MS) begin
                    key_state <= key_sync1; // ״̬ȷ��
                    cnt_debounce <= 0;
                end
            end else begin
                cnt_debounce <= 0;
            end
        end
    end

    // ===================== ���� / �̰���� =====================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cnt_hold  <= 32'd0;
            key_short <= 1'b0;
            key_long  <= 1'b0;
        end else begin
            // Ĭ���嵥��������
            key_short <= 1'b0;
            key_long  <= 1'b0;

            if (key_state == 1'b0) begin
                // �����ȶ������ڼ�
                if (cnt_hold < CNT_1S)
                    cnt_hold <= cnt_hold + 1;
                else
                    cnt_hold <= CNT_1S; // ����

                // ������ֵʱ�����������壨��һ�Σ�
                if (cnt_hold == CNT_1S - 1)
                    key_long <= 1'b1;
            end else begin
                // �ɿ�ʱ���������ʱ������ֵ���ڣ�������̰�����
                if ((cnt_hold > 0) && (cnt_hold < CNT_1S))
                    key_short <= 1'b1;

                // �ɿ����������
                cnt_hold <= 32'd0;
            end
        end
    end

endmodule